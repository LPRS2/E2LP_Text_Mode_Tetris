-----------------------------------------------------------------------------------
--  Odsek za racunarsku tehniku i medjuracunarske komunikacije                   --
--  Copyright � 2009 All Rights Reserved                                         --
--                                                                               --
--  Projekat: LabVezba2                                                          --
--  Ime modula: char_rom.vhd                                                     --
--  Autori: LPRS2 TIM 2009/2010 <LPRS2@KRT.neobee.net>                           --
--                                                                               --
--  Opis:                                                                        --
--          Char_rom generise tekst na ekranu.                                   --
--          Znak se predstavlja matricom 8x8 tacaka.                             --
--          Oblici znakova se nalaze u datoteci char_rom_def_mem.coe             --
--                                                                               --
-----------------------------------------------------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;



ENTITY char_rom IS PORT (
                         clk_i                : IN  STD_LOGIC;                            -- takt SIGNAL
                         character_address_i  : IN  STD_LOGIC_VECTOR (5 DOWNTO 0);        -- adresa karaktera
                         font_row_i           : IN  STD_LOGIC_VECTOR (2 DOWNTO 0);        -- ispis reda
                         font_col_i           : IN  STD_LOGIC_VECTOR (2 DOWNTO 0);        -- ispis kolone
                         rom_mux_output_o     : OUT STD_LOGIC                             -- izlazni SIGNAL iz char_rom-a
                        );
END char_rom;



ARCHITECTURE Behavioral OF char_rom IS

  SIGNAL rom_data    : STD_LOGIC_VECTOR( 7 DOWNTO 0 );       -- prosledjuje izlaz iz char_rom-a na ulaz u VGA
  SIGNAL rom_address : STD_LOGIC_VECTOR( 8 DOWNTO 0 );       -- preuzima character_address_i i font_row_i

	type t_mem is array(0 to 511) of std_logic_vector(7 downto 0);
	signal mem : t_mem := (
		"11111111",
		"10011001",
		"10011001",
		"11111111",
		"11111111",
		"10011001",
		"10011001",
		"11111111",
		"00011000",
		"00111100",
		"01100110",
		"01111110",
		"01100110",
		"01100110",
		"01100110",
		"00000000",
		"01111100",
		"01100110",
		"01100110",
		"01111100",
		"01100110",
		"01100110",
		"01111100",
		"00000000",
		"00111100",
		"01100110",
		"01100000",
		"01100000",
		"01100000",
		"01100110",
		"00111100",
		"00000000",
		"01111000",
		"01101100",
		"01100110",
		"01100110",
		"01100110",
		"01101100",
		"01111000",
		"00000000",
		"01111110",
		"01100000",
		"01100000",
		"01111000",
		"01100000",
		"01100000",
		"01111110",
		"00000000",
		"01111110",
		"01100000",
		"01100000",
		"01111000",
		"01100000",
		"01100000",
		"01100000",
		"00000000",
		"00111100",
		"01100110",
		"01100000",
		"01101110",
		"01100110",
		"01100110",
		"00111100",
		"00000000",
		"01100110",
		"01100110",
		"01100110",
		"01111110",
		"01100110",
		"01100110",
		"01100110",
		"00000000",
		"00111100",
		"00011000",
		"00011000",
		"00011000",
		"00011000",
		"00011000",
		"00111100",
		"00000000",
		"00011110",
		"00001100",
		"00001100",
		"00001100",
		"00001100",
		"01101100",
		"00111000",
		"00000000",
		"01100110",
		"01101100",
		"01111000",
		"01110000",
		"01111000",
		"01101100",
		"01100110",
		"00000000",
		"01100000",
		"01100000",
		"01100000",
		"01100000",
		"01100000",
		"01100000",
		"01111110",
		"00000000",
		"01100011",
		"01110111",
		"01111111",
		"01101011",
		"01100011",
		"01100011",
		"01100011",
		"00000000",
		"01100110",
		"01110110",
		"01111110",
		"01111110",
		"01101110",
		"01100110",
		"01100110",
		"00000000",
		"00111100",
		"01100110",
		"01100110",
		"01100110",
		"01100110",
		"01100110",
		"00111100",
		"00000000",
		"01111100",
		"01100110",
		"01100110",
		"01111100",
		"01100000",
		"01100000",
		"01100000",
		"00000000",
		"00111100",
		"01100110",
		"01100110",
		"01100110",
		"01100110",
		"00111100",
		"00001110",
		"00000000",
		"01111100",
		"01100110",
		"01100110",
		"01111100",
		"01111000",
		"01101100",
		"01100110",
		"00000000",
		"00111100",
		"01100110",
		"01100000",
		"00111100",
		"00000110",
		"01100110",
		"00111100",
		"00000000",
		"01111110",
		"00011000",
		"00011000",
		"00011000",
		"00011000",
		"00011000",
		"00011000",
		"00000000",
		"01100110",
		"01100110",
		"01100110",
		"01100110",
		"01100110",
		"01100110",
		"00111100",
		"00000000",
		"01100110",
		"01100110",
		"01100110",
		"01100110",
		"01100110",
		"00111100",
		"00011000",
		"00000000",
		"01100011",
		"01100011",
		"01100011",
		"01101011",
		"01111111",
		"01110111",
		"01100011",
		"00000000",
		"01100110",
		"01100110",
		"00111100",
		"00011000",
		"00111100",
		"01100110",
		"01100110",
		"00000000",
		"01100110",
		"01100110",
		"01100110",
		"00111100",
		"00011000",
		"00011000",
		"00011000",
		"00000000",
		"01111110",
		"00000110",
		"00001100",
		"00011000",
		"00110000",
		"01100000",
		"01111110",
		"00000000",
		"00111100",
		"00110000",
		"00110000",
		"00110000",
		"00110000",
		"00110000",
		"00111100",
		"00000000",
		"00011000",
		"00011000",
		"00011000",
		"00011000",
		"01111110",
		"00111100",
		"00011000",
		"00000000",
		"00111100",
		"00001100",
		"00001100",
		"00001100",
		"00001100",
		"00001100",
		"00111100",
		"00000000",
		"00000000",
		"00011000",
		"00111100",
		"01111110",
		"00011000",
		"00011000",
		"00011000",
		"00011000",
		"00000000",
		"00010000",
		"00110000",
		"01111111",
		"01111111",
		"00110000",
		"00010000",
		"00000000",
		"00000000",
		"00000000",
		"00000000",
		"00000000",
		"00000000",
		"00000000",
		"00000000",
		"00000000",
		"00011000",
		"00011000",
		"00011000",
		"00011000",
		"00000000",
		"00000000",
		"00011000",
		"00000000",
		"01100110",
		"01100110",
		"01100110",
		"00000000",
		"00000000",
		"00000000",
		"00000000",
		"00000000",
		"01100110",
		"01100110",
		"11111111",
		"01100110",
		"11111111",
		"01100110",
		"01100110",
		"00000000",
		"00011000",
		"00111110",
		"01100000",
		"00111100",
		"00000110",
		"01111100",
		"00011000",
		"00000000",
		"01100010",
		"01100110",
		"00001100",
		"00011000",
		"00110000",
		"01100110",
		"01000110",
		"00000000",
		"00111100",
		"01100110",
		"00111100",
		"00111000",
		"01100111",
		"01100110",
		"00111111",
		"00000000",
		"00000110",
		"00001100",
		"00011000",
		"00000000",
		"00000000",
		"00000000",
		"00000000",
		"00000000",
		"00001100",
		"00011000",
		"00110000",
		"00110000",
		"00110000",
		"00011000",
		"00001100",
		"00000000",
		"00110000",
		"00011000",
		"00001100",
		"00001100",
		"00001100",
		"00011000",
		"00110000",
		"00000000",
		"00000000",
		"01100110",
		"00111100",
		"11111111",
		"00111100",
		"01100110",
		"00000000",
		"00000000",
		"00000000",
		"00011000",
		"00011000",
		"01111110",
		"00011000",
		"00011000",
		"00000000",
		"00000000",
		"00000000",
		"00000000",
		"00000000",
		"00000000",
		"00000000",
		"00011000",
		"00011000",
		"00110000",
		"00000000",
		"00000000",
		"00000000",
		"01111110",
		"00000000",
		"00000000",
		"00000000",
		"00000000",
		"00000000",
		"00000000",
		"00000000",
		"00000000",
		"00000000",
		"00011000",
		"00011000",
		"00000000",
		"00000000",
		"00000011",
		"00000110",
		"00001100",
		"00011000",
		"00110000",
		"01100000",
		"00000000",
		"00111100",
		"01100110",
		"01101110",
		"01110110",
		"01100110",
		"01100110",
		"00111100",
		"00000000",
		"00011000",
		"00011000",
		"00111000",
		"00011000",
		"00011000",
		"00011000",
		"01111110",
		"00000000",
		"00111100",
		"01100110",
		"00000110",
		"00001100",
		"00110000",
		"01100000",
		"01111110",
		"00000000",
		"00111100",
		"01100110",
		"00000110",
		"00011100",
		"00000110",
		"01100110",
		"00111100",
		"00000000",
		"00000110",
		"00001110",
		"00011110",
		"01100110",
		"01111111",
		"00000110",
		"00000110",
		"00000000",
		"01111110",
		"01100000",
		"01111100",
		"00000110",
		"00000110",
		"01100110",
		"00111100",
		"00000000",
		"00111100",
		"01100110",
		"01100000",
		"01111100",
		"01100110",
		"01100110",
		"00111100",
		"00000000",
		"01111110",
		"01100110",
		"00001100",
		"00011000",
		"00011000",
		"00011000",
		"00011000",
		"00000000",
		"00111100",
		"01100110",
		"01100110",
		"00111100",
		"01100110",
		"01100110",
		"00111100",
		"00000000",
		"00111100",
		"01100110",
		"00111110",
		"00111110",
		"00000110",
		"01100110",
		"00111100",
		"00000000",
		"00011000",
		"00111100",
		"01100110",
		"01111110",
		"01100110",
		"01100110",
		"01100110",
		"00000000",
		"01111100",
		"01100110",
		"01100110",
		"01111100",
		"01100110",
		"01100110",
		"01111100",
		"00000000",
		"00111100",
		"01100110",
		"01100000",
		"01100000",
		"01100000",
		"01100110",
		"00111100",
		"00000000",
		"01111000",
		"01101100",
		"01100110",
		"01100110",
		"01100110",
		"01101100",
		"01111000",
		"00000000",
		"01111110",
		"01100000",
		"01100000",
		"01111110",
		"01100000",
		"01100000",
		"01111110",
		"00000000",
		"01111110",
		"01100000",
		"01100000",
		"01111000",
		"01100000",
		"01100000",
		"01100000",
		"00000000"
	);
	
	signal font_col_delayed: STD_LOGIC_VECTOR (2 DOWNTO 0);

BEGIN

                  ------------------|----------
                  --   ADDRESS      | OFFSET  |
                  ------------------|----------

	rom_address    <= character_address_i & font_row_i;

	process(clk_i)
	begin
		if rising_edge(clk_i) then
			rom_data <= mem(conv_integer(rom_address));
		end if;
	end process;

	process(clk_i)
	begin
		if rising_edge(clk_i) then
			font_col_delayed <= font_col_i;
		end if;
	end process;


PROCESS(font_col_delayed, rom_data) BEGIN

    CASE(font_col_delayed) IS

        WHEN  "000" => rom_mux_output_o <= rom_data(7);
        WHEN  "001" => rom_mux_output_o <= rom_data(6);
        WHEN  "010" => rom_mux_output_o <= rom_data(5);
        WHEN  "011" => rom_mux_output_o <= rom_data(4);
        WHEN  "100" => rom_mux_output_o <= rom_data(3);
        WHEN  "101" => rom_mux_output_o <= rom_data(2);
        WHEN  "110" => rom_mux_output_o <= rom_data(1);
        WHEN  "111" => rom_mux_output_o <= rom_data(0);
        WHEN OTHERS => rom_mux_output_o <= '0';

    END CASE;

END PROCESS;



END Behavioral;

